State|Population|Area
Alabama                   |4874747     |52420.07  
Alaska                    |739795       |665384.04
Arizona                   |7016270     |113990.30
Arkansas                  |3004279     |53178.55  
California                |39536653    |163696.32
Colorado                  |5607154     |104093.67
Connecticut               |3588184     |5543.41   
Delaware                  |961939       |2488.72   
Florida                   |20984400    |65757.70  
Georgia                   |10429379    |59425.15  
Hawaii                    |1427538     |10931.72  
Idaho                     |1716943     |83568.95  
Illinois                  |12802023    |57913.55  
Indiana                   |6666818     |36419.55  
Iowa                      |3145711     |56272.81  
Kansas                    |2913123     |82278.36  
Kentucky                  |4454189     |40407.80  
Louisiana                 |4684333     |52378.13  
Maine                     |1335907     |35379.74  
Maryland                  |6052177     |12405.93  
Massachusetts             |6859819     |10554.39  
Michigan                  |9962311     |96713.51
Minnesota                 |5576606     |86935.83  
Mississippi               |2984100     |48431.78  
Missouri                  |6113532     |69706.99  
Montana                   |1050493     |147039.71
Nebraska                  |1920076     |77347.81  
Nevada                    |2998039     |110571.82
New Hampshire             |1342795     |9349.16   
New Jersey                |9005644     |8722.58   
New Mexico                |2088070     |121590.30
New York                  |19849399    |54554.98  
North Carolina            |10273419    |53819.16  
North Dakota              |755393       |70698.32  
Ohio                      |11658609    |44825.58  
Oklahoma                  |3930864     |69898.87  
Oregon                    |4142776     |98378.54
Pennsylvania              |12805537    |46054.35  
Rhode Island              |1059639     |1544.89   
South Carolina            |5024369     |32020.49  
South Dakota              |869666       |77115.68  
Tennessee                 |6715984     |42144.25  
Texas                     |28304596    |268596.46
Utah                      |3101833     |84896.88  
Vermont                   |623657       |9616.36   
Virginia                  |8470020     |42774.93  
Washington                |7405743     |71297.95  
West Virginia             |1815857     |24230.04  
Wisconsin                 |5795483     |65496.38  
Wyoming                   |579315       |97813.01
